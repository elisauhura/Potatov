//  UART.v
//
//  Created by Elisa Silva on 26/10/21.
//  Copyright © 2021 Uhura. All rights reserved.

`include FIFO.v


// https://pbxbook.com/other/mac-tty.html


module UART_TX(
    reset,
    clock
);

endmodule

module UART_RX(
    rx,
    reset,
    clock
);

endmodule

module UART(
    cByte,
    cRead,
    cWrite,
    hByte,
    hCanRead,
    hCanWrite,
    tx,
    rx,
    reset,
    clock
);


endmodule
